module sbox(
    input inv,
    input [7:0] value,
    output reg [7:0] swap
);

always @(*)
    begin
        if (inv != 1)
            begin
                case (value)
                8'h00:swap <= 8'h63;
                8'h01:swap <= 8'h7c;
                8'h02:swap <= 8'h77;
                8'h03:swap <= 8'h7b;
                8'h04:swap <= 8'hf2;
                8'h05:swap <= 8'h6b;
                8'h06:swap <= 8'h6f;
                8'h07:swap <= 8'hc5;
                8'h08:swap <= 8'h30;
                8'h09:swap <= 8'h01;
                8'h0a:swap <= 8'h67;
                8'h0b:swap <= 8'h2b;
                8'h0c:swap <= 8'hfe;
                8'h0d:swap <= 8'hd7;
                8'h0e:swap <= 8'hab;
                8'h0f:swap <= 8'h76;
                8'h10:swap <= 8'hca;
                8'h11:swap <= 8'h82;
                8'h12:swap <= 8'hc9;
                8'h13:swap <= 8'h7d;
                8'h14:swap <= 8'hfa;
                8'h15:swap <= 8'h59;
                8'h16:swap <= 8'h47;
                8'h17:swap <= 8'hf0;
                8'h18:swap <= 8'had;
                8'h19:swap <= 8'hd4;
                8'h1a:swap <= 8'ha2;
                8'h1b:swap <= 8'haf;
                8'h1c:swap <= 8'h9c;
                8'h1d:swap <= 8'ha4;
                8'h1e:swap <= 8'h72;
                8'h1f:swap <= 8'hc0;
                8'h20:swap <= 8'hb7;
                8'h21:swap <= 8'hfd;
                8'h22:swap <= 8'h93;
                8'h23:swap <= 8'h26;
                8'h24:swap <= 8'h36;
                8'h25:swap <= 8'h3f;
                8'h26:swap <= 8'hf7;
                8'h27:swap <= 8'hcc;
                8'h28:swap <= 8'h34;
                8'h29:swap <= 8'ha5;
                8'h2a:swap <= 8'he5;
                8'h2b:swap <= 8'hf1;
                8'h2c:swap <= 8'h71;
                8'h2d:swap <= 8'hd8;
                8'h2e:swap <= 8'h31;
                8'h2f:swap <= 8'h15;
                8'h30:swap <= 8'h04;
                8'h31:swap <= 8'hc7;
                8'h32:swap <= 8'h23;
                8'h33:swap <= 8'hc3;
                8'h34:swap <= 8'h18;
                8'h35:swap <= 8'h96;
                8'h36:swap <= 8'h05;
                8'h37:swap <= 8'h9a;
                8'h38:swap <= 8'h07;
                8'h39:swap <= 8'h12;
                8'h3a:swap <= 8'h80;
                8'h3b:swap <= 8'he2;
                8'h3c:swap <= 8'heb;
                8'h3d:swap <= 8'h27;
                8'h3e:swap <= 8'hb2;
                8'h3f:swap <= 8'h75;
                8'h40:swap <= 8'h09;
                8'h41:swap <= 8'h83;
                8'h42:swap <= 8'h2c;
                8'h43:swap <= 8'h1a;
                8'h44:swap <= 8'h1b;
                8'h45:swap <= 8'h6e;
                8'h46:swap <= 8'h5a;
                8'h47:swap <= 8'ha0;
                8'h48:swap <= 8'h52;
                8'h49:swap <= 8'h3b;
                8'h4a:swap <= 8'hd6;
                8'h4b:swap <= 8'hb3;
                8'h4c:swap <= 8'h29;
                8'h4d:swap <= 8'he3;
                8'h4e:swap <= 8'h2f;
                8'h4f:swap <= 8'h84;
                8'h50:swap <= 8'h53;
                8'h51:swap <= 8'hd1;
                8'h52:swap <= 8'h00;
                8'h53:swap <= 8'hed;
                8'h54:swap <= 8'h20;
                8'h55:swap <= 8'hfc;
                8'h56:swap <= 8'hb1;
                8'h57:swap <= 8'h5b;
                8'h58:swap <= 8'h6a;
                8'h59:swap <= 8'hcb;
                8'h5a:swap <= 8'hbe;
                8'h5b:swap <= 8'h39;
                8'h5c:swap <= 8'h4a;
                8'h5d:swap <= 8'h4c;
                8'h5e:swap <= 8'h58;
                8'h5f:swap <= 8'hcf;
                8'h60:swap <= 8'hd0;
                8'h61:swap <= 8'hef;
                8'h62:swap <= 8'haa;
                8'h63:swap <= 8'hfb;
                8'h64:swap <= 8'h43;
                8'h65:swap <= 8'h4d;
                8'h66:swap <= 8'h33;
                8'h67:swap <= 8'h85;
                8'h68:swap <= 8'h45;
                8'h69:swap <= 8'hf9;
                8'h6a:swap <= 8'h02;
                8'h6b:swap <= 8'h7f;
                8'h6c:swap <= 8'h50;
                8'h6d:swap <= 8'h3c;
                8'h6e:swap <= 8'h9f;
                8'h6f:swap <= 8'ha8;
                8'h70:swap <= 8'h51;
                8'h71:swap <= 8'ha3;
                8'h72:swap <= 8'h40;
                8'h73:swap <= 8'h8f;
                8'h74:swap <= 8'h92;
                8'h75:swap <= 8'h9d;
                8'h76:swap <= 8'h38;
                8'h77:swap <= 8'hf5;
                8'h78:swap <= 8'hbc;
                8'h79:swap <= 8'hb6;
                8'h7a:swap <= 8'hda;
                8'h7b:swap <= 8'h21;
                8'h7c:swap <= 8'h10;
                8'h7d:swap <= 8'hff;
                8'h7e:swap <= 8'hf3;
                8'h7f:swap <= 8'hd2;
                8'h80:swap <= 8'hcd;
                8'h81:swap <= 8'h0c;
                8'h82:swap <= 8'h13;
                8'h83:swap <= 8'hec;
                8'h84:swap <= 8'h5f;
                8'h85:swap <= 8'h97;
                8'h86:swap <= 8'h44;
                8'h87:swap <= 8'h17;
                8'h88:swap <= 8'hc4;
                8'h89:swap <= 8'ha7;
                8'h8a:swap <= 8'h7e;
                8'h8b:swap <= 8'h3d;
                8'h8c:swap <= 8'h64;
                8'h8d:swap <= 8'h5d;
                8'h8e:swap <= 8'h19;
                8'h8f:swap <= 8'h73;
                8'h90:swap <= 8'h60;
                8'h91:swap <= 8'h81;
                8'h92:swap <= 8'h4f;
                8'h93:swap <= 8'hdc;
                8'h94:swap <= 8'h22;
                8'h95:swap <= 8'h2a;
                8'h96:swap <= 8'h90;
                8'h97:swap <= 8'h88;
                8'h98:swap <= 8'h46;
                8'h99:swap <= 8'hee;
                8'h9a:swap <= 8'hb8;
                8'h9b:swap <= 8'h14;
                8'h9c:swap <= 8'hde;
                8'h9d:swap <= 8'h5e;
                8'h9e:swap <= 8'h0b;
                8'h9f:swap <= 8'hdb;
                8'ha0:swap <= 8'he0;
                8'ha1:swap <= 8'h32;
                8'ha2:swap <= 8'h3a;
                8'ha3:swap <= 8'h0a;
                8'ha4:swap <= 8'h49;
                8'ha5:swap <= 8'h06;
                8'ha6:swap <= 8'h24;
                8'ha7:swap <= 8'h5c;
                8'ha8:swap <= 8'hc2;
                8'ha9:swap <= 8'hd3;
                8'haa:swap <= 8'hac;
                8'hab:swap <= 8'h62;
                8'hac:swap <= 8'h91;
                8'had:swap <= 8'h95;
                8'hae:swap <= 8'he4;
                8'haf:swap <= 8'h79;
                8'hb0:swap <= 8'he7;
                8'hb1:swap <= 8'hc8;
                8'hb2:swap <= 8'h37;
                8'hb3:swap <= 8'h6d;
                8'hb4:swap <= 8'h8d;
                8'hb5:swap <= 8'hd5;
                8'hb6:swap <= 8'h4e;
                8'hb7:swap <= 8'ha9;
                8'hb8:swap <= 8'h6c;
                8'hb9:swap <= 8'h56;
                8'hba:swap <= 8'hf4;
                8'hbb:swap <= 8'hea;
                8'hbc:swap <= 8'h65;
                8'hbd:swap <= 8'h7a;
                8'hbe:swap <= 8'hae;
                8'hbf:swap <= 8'h08;
                8'hc0:swap <= 8'hba;
                8'hc1:swap <= 8'h78;
                8'hc2:swap <= 8'h25;
                8'hc3:swap <= 8'h2e;
                8'hc4:swap <= 8'h1c;
                8'hc5:swap <= 8'ha6;
                8'hc6:swap <= 8'hb4;
                8'hc7:swap <= 8'hc6;
                8'hc8:swap <= 8'he8;
                8'hc9:swap <= 8'hdd;
                8'hca:swap <= 8'h74;
                8'hcb:swap <= 8'h1f;
                8'hcc:swap <= 8'h4b;
                8'hcd:swap <= 8'hbd;
                8'hce:swap <= 8'h8b;
                8'hcf:swap <= 8'h8a;
                8'hd0:swap <= 8'h70;
                8'hd1:swap <= 8'h3e;
                8'hd2:swap <= 8'hb5;
                8'hd3:swap <= 8'h66;
                8'hd4:swap <= 8'h48;
                8'hd5:swap <= 8'h03;
                8'hd6:swap <= 8'hf6;
                8'hd7:swap <= 8'h0e;
                8'hd8:swap <= 8'h61;
                8'hd9:swap <= 8'h35;
                8'hda:swap <= 8'h57;
                8'hdb:swap <= 8'hb9;
                8'hdc:swap <= 8'h86;
                8'hdd:swap <= 8'hc1;
                8'hde:swap <= 8'h1d;
                8'hdf:swap <= 8'h9e;
                8'he0:swap <= 8'he1;
                8'he1:swap <= 8'hf8;
                8'he2:swap <= 8'h98;
                8'he3:swap <= 8'h11;
                8'he4:swap <= 8'h69;
                8'he5:swap <= 8'hd9;
                8'he6:swap <= 8'h8e;
                8'he7:swap <= 8'h94;
                8'he8:swap <= 8'h9b;
                8'he9:swap <= 8'h1e;
                8'hea:swap <= 8'h87;
                8'heb:swap <= 8'he9;
                8'hec:swap <= 8'hce;
                8'hed:swap <= 8'h55;
                8'hee:swap <= 8'h28;
                8'hef:swap <= 8'hdf;
                8'hf0:swap <= 8'h8c;
                8'hf1:swap <= 8'ha1;
                8'hf2:swap <= 8'h89;
                8'hf3:swap <= 8'h0d;
                8'hf4:swap <= 8'hbf;
                8'hf5:swap <= 8'he6;
                8'hf6:swap <= 8'h42;
                8'hf7:swap <= 8'h68;
                8'hf8:swap <= 8'h41;
                8'hf9:swap <= 8'h99;
                8'hfa:swap <= 8'h2d;
                8'hfb:swap <= 8'h0f;
                8'hfc:swap <= 8'hb0;
                8'hfd:swap <= 8'h54;
                8'hfe:swap <= 8'hbb;
                8'hff:swap <= 8'h16;
                default: 
                swap = 0;
            endcase
            end
    else
        begin
            case (value)
                8'h00:swap <= 8'h52;
                8'h01:swap <= 8'h09;
                8'h02:swap <= 8'h6a;
                8'h03:swap <= 8'hd5;
                8'h04:swap <= 8'h30;
                8'h05:swap <= 8'h36;
                8'h06:swap <= 8'ha5;
                8'h07:swap <= 8'h38;
                8'h08:swap <= 8'hbf;
                8'h09:swap <= 8'h40;
                8'h0a:swap <= 8'ha3;
                8'h0b:swap <= 8'h9e;
                8'h0c:swap <= 8'h81;
                8'h0d:swap <= 8'hf3;
                8'h0e:swap <= 8'hd7;
                8'h0f:swap <= 8'hfb;
                8'h10:swap <= 8'h7c;
                8'h11:swap <= 8'he3;
                8'h12:swap <= 8'h39;
                8'h13:swap <= 8'h82;
                8'h14:swap <= 8'h9b;
                8'h15:swap <= 8'h2f;
                8'h16:swap <= 8'hff;
                8'h17:swap <= 8'h87;
                8'h18:swap <= 8'h34;
                8'h19:swap <= 8'h8e;
                8'h1a:swap <= 8'h43;
                8'h1b:swap <= 8'h44;
                8'h1c:swap <= 8'hc4;
                8'h1d:swap <= 8'hde;
                8'h1e:swap <= 8'he9;
                8'h1f:swap <= 8'hcb;
                8'h20:swap <= 8'h54;
                8'h21:swap <= 8'h7b;
                8'h22:swap <= 8'h94;
                8'h23:swap <= 8'h32;
                8'h24:swap <= 8'ha6;
                8'h25:swap <= 8'hc2;
                8'h26:swap <= 8'h23;
                8'h27:swap <= 8'h3d;
                8'h28:swap <= 8'hee;
                8'h29:swap <= 8'h4c;
                8'h2a:swap <= 8'h95;
                8'h2b:swap <= 8'h0b;
                8'h2c:swap <= 8'h42;
                8'h2d:swap <= 8'hfa;
                8'h2e:swap <= 8'hc3;
                8'h2f:swap <= 8'h4e;
                8'h30:swap <= 8'h08;
                8'h31:swap <= 8'h2e;
                8'h32:swap <= 8'ha1;
                8'h33:swap <= 8'h66;
                8'h34:swap <= 8'h28;
                8'h35:swap <= 8'hd9;
                8'h36:swap <= 8'h24;
                8'h37:swap <= 8'hb2;
                8'h38:swap <= 8'h76;
                8'h39:swap <= 8'h5b;
                8'h3a:swap <= 8'ha2;
                8'h3b:swap <= 8'h49;
                8'h3c:swap <= 8'h6d;
                8'h3d:swap <= 8'h8b;
                8'h3e:swap <= 8'hd1;
                8'h3f:swap <= 8'h25;
                8'h40:swap <= 8'h72;
                8'h41:swap <= 8'hf8;
                8'h42:swap <= 8'hf6;
                8'h43:swap <= 8'h64;
                8'h44:swap <= 8'h86;
                8'h45:swap <= 8'h68;
                8'h46:swap <= 8'h98;
                8'h47:swap <= 8'h16;
                8'h48:swap <= 8'hd4;
                8'h49:swap <= 8'ha4;
                8'h4a:swap <= 8'h5c;
                8'h4b:swap <= 8'hcc;
                8'h4c:swap <= 8'h5d;
                8'h4d:swap <= 8'h65;
                8'h4e:swap <= 8'hb6;
                8'h4f:swap <= 8'h92;
                8'h50:swap <= 8'h6c;
                8'h51:swap <= 8'h70;
                8'h52:swap <= 8'h48;
                8'h53:swap <= 8'h50;
                8'h54:swap <= 8'hfd;
                8'h55:swap <= 8'hed;
                8'h56:swap <= 8'hb9;
                8'h57:swap <= 8'hda;
                8'h58:swap <= 8'h5e;
                8'h59:swap <= 8'h15;
                8'h5a:swap <= 8'h46;
                8'h5b:swap <= 8'h57;
                8'h5c:swap <= 8'ha7;
                8'h5d:swap <= 8'h8d;
                8'h5e:swap <= 8'h9d;
                8'h5f:swap <= 8'h84;
                8'h60:swap <= 8'h90;
                8'h61:swap <= 8'hd8;
                8'h62:swap <= 8'hab;
                8'h63:swap <= 8'h00;
                8'h64:swap <= 8'h8c;
                8'h65:swap <= 8'hbc;
                8'h66:swap <= 8'hd3;
                8'h67:swap <= 8'h0a;
                8'h68:swap <= 8'hf7;
                8'h69:swap <= 8'he4;
                8'h6a:swap <= 8'h58;
                8'h6b:swap <= 8'h05;
                8'h6c:swap <= 8'hb8;
                8'h6d:swap <= 8'hb3;
                8'h6e:swap <= 8'h45;
                8'h6f:swap <= 8'h06;
                8'h70:swap <= 8'hd0;
                8'h71:swap <= 8'h2c;
                8'h72:swap <= 8'h1e;
                8'h73:swap <= 8'h8f;
                8'h74:swap <= 8'hca;
                8'h75:swap <= 8'h3f;
                8'h76:swap <= 8'h0f;
                8'h77:swap <= 8'h02;
                8'h78:swap <= 8'hc1;
                8'h79:swap <= 8'haf;
                8'h7a:swap <= 8'hbd;
                8'h7b:swap <= 8'h03;
                8'h7c:swap <= 8'h01;
                8'h7d:swap <= 8'h13;
                8'h7e:swap <= 8'h8a;
                8'h7f:swap <= 8'h6b;
                8'h80:swap <= 8'h3a;
                8'h81:swap <= 8'h91;
                8'h82:swap <= 8'h11;
                8'h83:swap <= 8'h41;
                8'h84:swap <= 8'h4f;
                8'h85:swap <= 8'h67;
                8'h86:swap <= 8'hdc;
                8'h87:swap <= 8'hea;
                8'h88:swap <= 8'h97;
                8'h89:swap <= 8'hf2;
                8'h8a:swap <= 8'hcf;
                8'h8b:swap <= 8'hce;
                8'h8c:swap <= 8'hf0;
                8'h8d:swap <= 8'hb4;
                8'h8e:swap <= 8'he6;
                8'h8f:swap <= 8'h73;
                8'h90:swap <= 8'h96;
                8'h91:swap <= 8'hac;
                8'h92:swap <= 8'h74;
                8'h93:swap <= 8'h22;
                8'h94:swap <= 8'he7;
                8'h95:swap <= 8'had;
                8'h96:swap <= 8'h35;
                8'h97:swap <= 8'h85;
                8'h98:swap <= 8'he2;
                8'h99:swap <= 8'hf9;
                8'h9a:swap <= 8'h37;
                8'h9b:swap <= 8'he8;
                8'h9c:swap <= 8'h1c;
                8'h9d:swap <= 8'h75;
                8'h9e:swap <= 8'hdf;
                8'h9f:swap <= 8'h6e;
                8'ha0:swap <= 8'h47;
                8'ha1:swap <= 8'hf1;
                8'ha2:swap <= 8'h1a;
                8'ha3:swap <= 8'h71;
                8'ha4:swap <= 8'h1d;
                8'ha5:swap <= 8'h29;
                8'ha6:swap <= 8'hc5;
                8'ha7:swap <= 8'h89;
                8'ha8:swap <= 8'h6f;
                8'ha9:swap <= 8'hb7;
                8'haa:swap <= 8'h62;
                8'hab:swap <= 8'h0e;
                8'hac:swap <= 8'haa;
                8'had:swap <= 8'h18;
                8'hae:swap <= 8'hbe;
                8'haf:swap <= 8'h1b;
                8'hb0:swap <= 8'hfc;
                8'hb1:swap <= 8'h56;
                8'hb2:swap <= 8'h3e;
                8'hb3:swap <= 8'h4b;
                8'hb4:swap <= 8'hc6;
                8'hb5:swap <= 8'hd2;
                8'hb6:swap <= 8'h79;
                8'hb7:swap <= 8'h20;
                8'hb8:swap <= 8'h9a;
                8'hb9:swap <= 8'hdb;
                8'hba:swap <= 8'hc0;
                8'hbb:swap <= 8'hfe;
                8'hbc:swap <= 8'h78;
                8'hbd:swap <= 8'hcd;
                8'hbe:swap <= 8'h5a;
                8'hbf:swap <= 8'hf4;
                8'hc0:swap <= 8'h1f;
                8'hc1:swap <= 8'hdd;
                8'hc2:swap <= 8'ha8;
                8'hc3:swap <= 8'h33;
                8'hc4:swap <= 8'h88;
                8'hc5:swap <= 8'h07;
                8'hc6:swap <= 8'hc7;
                8'hc7:swap <= 8'h31;
                8'hc8:swap <= 8'hb1;
                8'hc9:swap <= 8'h12;
                8'hca:swap <= 8'h10;
                8'hcb:swap <= 8'h59;
                8'hcc:swap <= 8'h27;
                8'hcd:swap <= 8'h80;
                8'hce:swap <= 8'hec;
                8'hcf:swap <= 8'h5f;
                8'hd0:swap <= 8'h60;
                8'hd1:swap <= 8'h51;
                8'hd2:swap <= 8'h7f;
                8'hd3:swap <= 8'ha9;
                8'hd4:swap <= 8'h19;
                8'hd5:swap <= 8'hb5;
                8'hd6:swap <= 8'h4a;
                8'hd7:swap <= 8'h0d;
                8'hd8:swap <= 8'h2d;
                8'hd9:swap <= 8'he5;
                8'hda:swap <= 8'h7a;
                8'hdb:swap <= 8'h9f;
                8'hdc:swap <= 8'h93;
                8'hdd:swap <= 8'hc9;
                8'hde:swap <= 8'h9c;
                8'hdf:swap <= 8'hef;
                8'he0:swap <= 8'ha0;
                8'he1:swap <= 8'he0;
                8'he2:swap <= 8'h3b;
                8'he3:swap <= 8'h4d;
                8'he4:swap <= 8'hae;
                8'he5:swap <= 8'h2a;
                8'he6:swap <= 8'hf5;
                8'he7:swap <= 8'hb0;
                8'he8:swap <= 8'hc8;
                8'he9:swap <= 8'heb;
                8'hea:swap <= 8'hbb;
                8'heb:swap <= 8'h3c;
                8'hec:swap <= 8'h83;
                8'hed:swap <= 8'h53;
                8'hee:swap <= 8'h99;
                8'hef:swap <= 8'h61;
                8'hf0:swap <= 8'h17;
                8'hf1:swap <= 8'h2b;
                8'hf2:swap <= 8'h04;
                8'hf3:swap <= 8'h7e;
                8'hf4:swap <= 8'hba;
                8'hf5:swap <= 8'h77;
                8'hf6:swap <= 8'hd6;
                8'hf7:swap <= 8'h26;
                8'hf8:swap <= 8'he1;
                8'hf9:swap <= 8'h69;
                8'hfa:swap <= 8'h14;
                8'hfb:swap <= 8'h63;
                8'hfc:swap <= 8'h55;
                8'hfd:swap <= 8'h21;
                8'hfe:swap <= 8'h0c;
                8'hff:swap <= 8'h7d;
                default: 
                swap = 0;
            endcase
        end
    end


endmodule