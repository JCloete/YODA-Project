module uVader(
    input clk,
    input reset,
    input  start,
    output reg [2:0]led, //RGB led (to be linked state in HW)
    output reg [2:0]state
);

// key = [113, 113, 113, 113, 119, 119, 119, 119, 101, 101, 101, 101, 114, 114, 116, 121]
// arr = [68, 105, 115, 99, 111, 109, 98, 111, 98, 117, 108, 97, 116, 101, 109, 101]
    reg [7:0] arr [15:0]; // The array with the data
    reg [7:0] key [15:0]; // The array with the key
    reg invert = 1;
    reg [7:0] in;
    wire [7:0] out;
    integer d = 0;
    
    // ----------          ----- FUNCTION DECLARATIONS -----         ----------//
    sbox mut(clk,invert, in, out);
    
    function addKey;
        input inv;
        integer i;
        begin
            i = 0;
            while (i < 128) begin
                arr[i] = arr[i] ^ key[i];
                i = i + 1;
            end
        end
    endfunction
    
    function subBytes;
        input inv;
        input incoming_byte;
        begin
            in = incoming_byte;
            subBytes = out;
        end
    endfunction

    function shiftRows;
        input inv;
        integer f,j,t;
        integer c;
        begin
            c = 1;
            for (f = 0; f < 4; f = f + 1)
                begin
                    if (inv == 0) begin
                        while (c < f) begin
                            t = arr[f*4];
                            arr[(f*4) + 0] = arr[(f*4) + 1]; arr[(f*4) + 1] = arr[(f*4) + 2]; arr[(f*4) + 2] = arr[(f*4) + 3]; arr[(f*4) + 3] = t;
                            c = c + 1;
                        end
                        c = 0;
                    end else begin
                        for (j = 0;j < 3 ;j = j + 1 ) begin
                            while (c < f) begin
                            t = arr[f*4];
                            arr[(f*4) + 0] = arr[(f*4) + 1]; arr[(f*4) + 1] = arr[(f*4) + 2]; arr[(f*4) + 2] = arr[(f*4) + 3]; arr[(f*4) + 3] = t;
                            c = c + 1;
                        end
                        c = 0;
                        end
                    end
                end
        end
    endfunction
    
    function [7:0]galois;
        input[7:0] a;
        input[7:0] b;
        reg[7:0] p;
        reg[7:0] highBit;
        begin
            p = 0;
            highBit = 0;
            repeat (8) begin
                if ((b & 1) == 1) begin
                    p = p ^ a;
                end
                highBit = a & 8'h80;
                a = a << 1;
                if (highBit == 8'h80) begin
                    a = a ^ 8'h1b;
                end
                b = b >> 1;
            end
            galois = p % 256;
        end
    endfunction

    function mixColumns;
        input inv;
        reg [7:0] temp [3:0];
        integer count;
        reg [3:0] a,b,c,d;
        begin
            if (inv == 0) begin
                for (count = 0; count < 4; count = count + 1) begin
                    a = count + 0; b = count + 4; c = count + 8; d = count + 12;
                    temp[0] = arr[a]; temp[1] = arr[b]; temp[2] = arr[c]; temp[3] = arr[d];
                    arr[a] = galois(temp[0], 2) ^ galois(temp[3], 1) ^ galois(temp[2], 1) ^ galois(temp[1], 3);
                    arr[b] = galois(temp[1], 2) ^ galois(temp[0], 1) ^ galois(temp[3], 1) ^ galois(temp[2], 3);
                    arr[c] = galois(temp[2], 2) ^ galois(temp[1], 1) ^ galois(temp[0], 1) ^ galois(temp[3], 3);
                    arr[d] = galois(temp[3], 2) ^ galois(temp[2], 1) ^ galois(temp[1], 1) ^ galois(temp[0], 3);
                end
            end else begin
                for (count = 0; count < 4; count = count + 1) begin
                    a = count + 0; b = count + 4; c = count + 8; d = count + 12;
                    temp[0] = arr[a]; temp[1] = arr[b]; temp[2] = arr[c]; temp[3] = arr[d];
                    arr[a] = galois(temp[0], 14) ^ galois(temp[3], 9) ^ galois(temp[2], 13) ^ galois(temp[1], 11);
                    arr[b] = galois(temp[1], 14) ^ galois(temp[0], 9) ^ galois(temp[3], 13) ^ galois(temp[2], 11);
                    arr[c] = galois(temp[2], 14) ^ galois(temp[1], 9) ^ galois(temp[0], 13) ^ galois(temp[3], 11);
                    arr[d] = galois(temp[3], 14) ^ galois(temp[2], 9) ^ galois(temp[1], 13) ^ galois(temp[0], 11);
            end
            end
        end
    endfunction

    function round;
        input inv;
        integer dump, i;
        begin
            if (inv == 1) begin
                dump = addKey(inv);
                dump = mixColumns(inv);
                dump = shiftRows(inv);
                for (i=0; i < 16; i = i + 1) begin
                    dump = subBytes(inv, arr[i]);
                end
            end
            else begin
                for (i=0; i < 16; i = i + 1) begin
                    dump = subBytes(inv, arr[i]);
                end
                dump = shiftRows(inv);
                dump = mixColumns(inv);
                dump = addKey(inv);
            end
        end 
    endfunction

    function crypt; // 1 will decrypt, 0 will encrypt
        input inv;
        integer r,i,dump;
        begin
            if (inv == 1) begin
                dump = addKey(inv);
                dump = shiftRows(inv);
                for (i=0; i < 16; i = i + 1) begin
                    dump = subBytes(inv, arr[i]);
                end
                for (r = 0; r < 9; r = r+1) begin
                    dump = round(inv);
                end
                dump = addKey(inv);
            end
            else begin
                dump = addKey(inv);
                for (r = 0; r < 9; r = r+1) begin
                    dump = round(inv);
                end
                for (i=0; i < 16; i = i + 1) begin
                    dump = subBytes(inv, arr[i]);
                end
                dump = shiftRows(inv);
                dump = addKey(inv);
            end
        end
        
    endfunction

    always @(posedge reset) begin
        arr[0] = 204;
        arr[1] = 110;
        arr[2] = 219;
        arr[3] = 177;
        arr[4] = 21;
        arr[5] = 152;
        arr[6] = 49;
        arr[7] = 113;
        arr[8] = 39;
        arr[9] = 162;
        arr[10] = 150;
        arr[11] = 37;
        arr[12] = 144;
        arr[13] = 24;
        arr[14] = 51;
        arr[15] = 210;
        key[0] = 113;
        key[1] = 113;
        key[2] = 113;
        key[3] = 113;
        key[4] = 119;
        key[5] = 119;
        key[6] = 119;
        key[7] = 119;
        key[8] = 101;
        key[9] = 101;
        key[10] = 101;
        key[11] = 101;
        key[12] = 114;
        key[13] = 114;
        key[14] = 116;
        key[15] = 121;
    end

    integer i;
    always @(posedge start) begin
        // d = crypt(1);
        $display("Start Array");
        for (i = 0; i < 16; i = i + 4)
            begin
                $display("%3d %3d %3d %3d",arr[i], arr[i + 1], arr[i + 2], arr[i + 3]);
            end
        
        $display("\nAdd Key");
        d = addKey(1);
        for (i = 0; i < 16; i = i + 4)
            begin
                $display("%3d %3d %3d %3d",arr[i], arr[i + 1], arr[i + 2], arr[i + 3]);
            end

        $display("\nShift Rows");
        d = shiftRows(1);
        for (i = 0; i < 16; i = i + 4)
            begin
                $display("%3d %3d %3d %3d",arr[i], arr[i + 1], arr[i + 2], arr[i + 3]);
            end

        $display("\nSub Bytes");
        for (i=0; i < 16; i = i + 1) begin
                d = subBytes(1, arr[i]);
            end
        for (i = 0; i < 16; i = i + 4)
            begin
                $display("%3d %3d %3d %3d",arr[i], arr[i + 1], arr[i + 2], arr[i + 3]);
            end
        
        $display("\nMix Columns");
        d = mixColumns(1);
        for (i = 0; i < 16; i = i + 4)
            begin
                $display("%3d %3d %3d %3d",arr[i], arr[i + 1], arr[i + 2], arr[i + 3]);
            end
        
        
        // d = crypt(0);
        // $display("\n-- Start array --\n");
        // for (i = 0; i < 16; i = i + 4)
        //     begin
        //         $display("%3d %3d %3d %3d",arr[i], arr[i + 1], arr[i + 2], arr[i + 3]);
        //     end
        // if crypt(1) we expect:
        // 68 105 115  99
        // 111 109  98 111
        // 98 117 108  97
        // 116 101 109 101
    end
    // ----------          ----- ----    -----    ---- -----         ----------//
endmodule // 