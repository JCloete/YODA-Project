module SD_SIM(
    input clka,
    input ena,
    input [0 : 0] wea,
    input [3 : 0] addra,
    input [127 : 0] dina,
    output reg [127 : 0] douta
);

reg [127:0] source [8:0];

initial begin
    source[0] = 11001100011011101101101110110001000101011001100000110001011100010010011110100010100101100010010110010000000110000011001111010010;
    source[1] = 01110001011100010111000101110001011101110111011101110111011101110110010101100101011001010110010101110010011100100111010001111001;
    source[2] = 01110001011100010111000101110001011101110111011101110111011101110110010101100101011001010110010101110010011100100111010001111001;
    source[3] = 01101011011001010111100101100010011011110110000101110010011001000111011101100001011100100111001001101001011011110111001001110011;
    source[4] = 01010011011101000111010101110000011001010110111001100100011011110111010101110011011101000111001001100101011001010111001100110101;
    source[5] = 01010100011010000110010101010111011010010110111001100010011001010111001001100111011101010110110001100001011100100111001100110010;
    source[6] = 01000100011010010111001101100011011011110110110101100010011011110110001001110101011011000110000101110100011001010110110101100101;
    source[7] = 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end

always @(posedge clka) begin
    if (wea) begin
        source[addra] <= dina;
    end else begin
        douta <= source[addra];
    end
end

endmodule